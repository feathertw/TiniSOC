// tag:20 index:6 offset:4 word:2
`define TAG  20
`define IDX   6
`define OFS   4
`define BLK 512
`define DEP  64
`define WOR  32
`include "ram_tag.v"
`include "ram_valid.v"
`include "ram_data.v"

module icache(
);
endmodule

